signature sGreet { ER greetInKlingon(void); };

// Generate an RPC client proxy for the signature. The output looks like the
// following:
//
//     composite tGreetClientProxy {
//         entry sGreet eEntry;
//         call sChannel cChannel;
//         /* ... */
//     }
//
//     composite tGreetServerProxy {
//         call sGreet cEntry;
//         call sChannel cChannel;
//         entry sUnmarshalerMain  eService;
//         /* ... */
//     }
//
generate(AbstractRPCProxyPlugin, sGreet,
         "clientCelltypeName = tGreetClientProxy, "
         "serverCelltypeName = tGreetServerProxy, ");

// Import the definitions of kernel objects
import(<kernel.cdl>);

// System services
import("syssvc/tSerialPort.cdl");
import("syssvc/tSysLog.cdl");
import("syssvc/tSysLogAdapter.cdl");
import("syssvc/tLogTask.cdl");
import("syssvc/tBanner.cdl");

// Target-specific part
import("target.cdl");

//////////////////////////////////////////////////////////////////////////
//
// Syslog facility
//
//////////////////////////////////////////////////////////////////////////

cell tSysLogAdapter SysLogAdapter {
    cSysLog = rKernelDomain::SysLog.eSysLog;
};

region rKernelDomain {

cell tSysLog SysLog {
    logBufferSize = 32;                 /* ログバッファのサイズ */
    initLogMask = C_EXP("LOG_UPTO(LOG_NOTICE)");
                                        /* ログバッファに記録すべき重要度 */
    initLowMask = C_EXP("LOG_UPTO(LOG_EMERG)");
                                        /* 低レベル出力すべき重要度 */
    /* 低レベル出力との結合 */
    cPutLog = PutLogTarget.ePutLog;
};

[restrict(eSerialPort={rKernelDomain})]
cell tSerialPort SerialPort1 {
    receiveBufferSize = 256;            /* 受信バッファのサイズ */
    sendBufferSize    = 256;            /* 送信バッファのサイズ */

    /* ターゲット依存部との結合 */
    cSIOPort = SIOPortTarget1.eSIOPort;
    eiSIOCBR <= SIOPortTarget1.ciSIOCBR;    /* コールバック */
};

cell tLogTask LogTask {
    priority  = 3;                  /* システムログタスクの優先度 */
    stackSize = LogTaskStackSize;   /* システムログタスクのスタックサイズ */

    /* シリアルインタフェースドライバとの結合 */
    cSerialPort        = SerialPort1.eSerialPort;
    cnSerialPortManage = SerialPort1.enSerialPortManage;

    /* システムログ機能との結合 */
    cSysLog = SysLog.eSysLog;

    /* 低レベル出力との結合 */
    cPutLog = PutLogTarget.ePutLog;
};

cell tBanner Banner {
    /* 属性の設定 */
    targetName      = BannerTargetName;
    copyrightNotice = BannerCopyrightNotice;
};

}; // region rKernelDomain

//////////////////////////////////////////////////////////////////////////
//
// Main application
//
//////////////////////////////////////////////////////////////////////////

[singleton]
celltype tApp {
    require tKernel.eKernel;

    /// The entry point
    entry sTaskBody eMain;
};

cell tKernel HRPKernel {};

cell tApp App {};

[domain(HRP, "user")]
region rAppDomain {

cell tTask MainTask {
    cTaskBody = App.eMain;
    attribute = C_EXP("TA_ACT");
    priority = C_EXP("MAIN_PRIORITY");
    stackSize = C_EXP("STACK_SIZE");
};

}; // region rAppDomain
